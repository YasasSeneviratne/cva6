module rm_tb_top #(
	parameter NUM_EVENTS	= 4,
	parameter NUM_LANES	= 4,
	parameter NUM_RULES	= 5
	)(
	input 				clk_i,
	input 				rst_ni_tb,
	input [NUM_EVENTS-1:0]		signal_tb, //random event signal
	input [NUM_EVENTS-1:0]		reset_lane_i_tb,
//	output ariane_pkg::lane_ctrl 		lane_cnt_o,
//	input ariane_pkg::runtime_monitor_ctrl	[NUM_EVENTS-1:0] rm_cnt_i,
	input [riscv::VLEN-1:0]	    	pc_i_tb,
	input  				enque_ins_tb,
	input [6:0]			opcode_i_tb,

//	output logic [NUM_EVENTS-1:0][NUM_LANES-1:0]	lane_vector,
//	output logic [NUM_LANES-1:0]			lane_reset
	output logic [NUM_EVENTS-1:0]	lane_vector_0,
	output logic [NUM_EVENTS-1:0]	lane_vector_1,
	output logic [NUM_EVENTS-1:0]	lane_vector_2,
	output logic [NUM_EVENTS-1:0]	lane_vector_3,
	
	output logic [NUM_RULES-1:0]	monitor_o_0,
	output logic [NUM_RULES-1:0]	monitor_o_1,
	output logic [NUM_RULES-1:0]	monitor_o_2,
	output logic [NUM_RULES-1:0]	monitor_o_3,
	
	output logic [NUM_LANES-1:0]   lane_reset,
	output logic [NUM_LANES-1:0]   lane_reset_0,
	output logic [NUM_LANES-1:0]   lane_reset_1,
	output logic [NUM_LANES-1:0]   lane_reset_2,
	output logic [NUM_LANES-1:0]   lane_reset_3
	);

	ariane_pkg::lane_ctrl [NUM_EVENTS-1: 0]        rm_event_o;

	ariane_pkg::runtime_monitor_ctrl	[NUM_EVENTS-1:0] rm_cnt;
	ariane_pkg::runtime_monitor_ctrl	rm_cnt_o;

	logic [NUM_LANES-1: 0][NUM_RULES-1:0]	monitor_o;
	logic [NUM_EVENTS-1:0][NUM_LANES-1:0]	lane_vector;
	//logic [NUM_LANES-1:0]			lane_reset;


	//--------- SIMULATION SUPPORT---------------
	//Indexing not supported in verilator :(
	assign lane_vector_0 = lane_vector[0];
	assign lane_vector_1 = lane_vector[1];
	assign lane_vector_2 = lane_vector[2];
	assign lane_vector_3 = lane_vector[3];

	assign monitor_o_0 = monitor_o[0];
	assign monitor_o_1 = monitor_o[1];
	assign monitor_o_2 = monitor_o[2];
	assign monitor_o_3 = monitor_o[3];

	assign lane_reset_0 = lane_reset[0];	
	assign lane_reset_1 = lane_reset[1];	
	assign lane_reset_2 = lane_reset[2];	
	assign lane_reset_3 = lane_reset[3];	
	//Input sygnals must be sunchronoized to observe correct behaviour

	logic				rst_ni;
	logic [NUM_EVENTS-1:0]		signal;
	logic [NUM_EVENTS-1:0]		reset_lane_i;
	logic [riscv::VLEN-1:0]    	pc_i;
	logic 				enque_ins;
	logic [6:0]			opcode_i;

	always_ff @(posedge clk_i) begin
		rst_ni		<= rst_ni_tb;
		signal		<= signal_tb;
		reset_lane_i	<= reset_lane_i_tb;
		pc_i 		<= pc_i_tb;
		enque_ins	<= enque_ins_tb;
		opcode_i	<= opcode_i_tb;
	end
	/////////////////////////////////////////////////
	
	always_ff @(posedge clk_i , negedge rst_ni) begin
		if (!rst_ni) begin
			rm_cnt <= '0;
		end 
		else begin
			for (int i=0; i<NUM_EVENTS-1; i++) begin
				rm_cnt[i+1] <= rm_cnt[i];
			end
			rm_cnt[0] <= rm_cnt_o;
		        //in cof1 number of lanes == events therfore	
                        for (int i=0; i<NUM_EVENTS; i++) begin
                                if(reset_lane_i[i])
				     rm_cnt[i+1] <= '0;
			end
		end		
	end


	genvar i;
	generate
		for(i=0; i<NUM_EVENTS-1; i++) begin
			rm_event_detector #(
			.NUM_VARS(1),
			.NUM_LANES
			)
			ev (
			.clk_i,
			.rst_ni,
			.signal(signal[i]),
			.ref_val(1'b1),
			.rm_cnt_i(rm_cnt[i]),
			.lane_cnt_o(rm_event_o[i]),
			.reset_lane_i(reset_lane_i[i])
			);	
		end
	endgenerate
	

	//rm_event_detector #(
	//.NUM_VARS(1),
	//.NUM_LANES
	//)
	//ev1 (
	//.signal(signal[1]),
	//.ref_val(1'b1),
	//.rm_cnt_i(rm_cnt[1]),
	//.lane_cnt_o(rm_event_o[1]),
	//.reset_lane_i(reset_lane_i[1])
	//);	
	
	rm_event_detector #(
	.NUM_VARS(1),
	.NUM_LANES,
	.LEAF_EVENT(1)
	)
	ev (
	.clk_i,
	.rst_ni,
	.signal(signal[NUM_EVENTS-1]),
	.ref_val(1'b1),
	.rm_cnt_i(rm_cnt[NUM_EVENTS-1]),
	.lane_cnt_o(rm_event_o[NUM_EVENTS-1]),
	.reset_lane_i(reset_lane_i[NUM_EVENTS-1])
	);	


	rm_lane_allocator #(
	.NUM_LANES,
	.NUM_EVENTS
	)
	rm_alloc (
	.clk_i,
	.rst_ni,
	.flush_i(0),
	.opcode	(opcode_i),
	.pc_i,
	.reset_monitor (rm_event_o),
	.entry_queued_i (enque_ins),
	.monitor_o (rm_cnt_o)
	);


	rm_event_router #(
	.NUM_LANES,
	.NUM_EVENTS
	)
	router (
	.events_i	(rm_event_o),
	.lane_vector_o (lane_vector),
	.lane_reset_o (lane_reset)
	);
	
	rm_monitor  #(
	.NUM_LANES,
	.NUM_EVENTS, 
	.NUM_RULES
	)	
	rm(
	.clk_i,
	.rst_ni,
	.lane_vector_i(lane_vector),
	.lane_reset_i(lane_reset),
	.monitor_o
	);
	

endmodule
