




/*
******************** Summary ********************
report for ltl0c0
Number of nodes = 9
Number of edges = 17
Average edge per node = 0.529411764706
Number of start nodes = 3
Number of report nodes = 4
does have all_input = False
does have special element = False
is Homogenous = True
stride value = 1
Max Fan-in = 4
Max Fan-out = 3
Max value in dim = 255
average number of intervals per STE = 2.11111111111
#######################################################
*/

 



module LUT_Match_ltl0c0_1 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd0) &&(input_capture[7:0] <= 8'd1) && 1'b1) ||
     ((input_capture[7:0] >= 8'd8) &&(input_capture[7:0] <= 8'd9) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_2 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd2) &&(input_capture[7:0] <= 8'd3) && 1'b1) ||
     ((input_capture[7:0] >= 8'd6) &&(input_capture[7:0] <= 8'd7) && 1'b1) ||
     ((input_capture[7:0] >= 8'd10) &&(input_capture[7:0] <= 8'd11) && 1'b1) ||
     ((input_capture[7:0] >= 8'd14) &&(input_capture[7:0] <= 8'd15) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_3 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd4) &&(input_capture[7:0] <= 8'd5) && 1'b1) ||
     ((input_capture[7:0] >= 8'd12) &&(input_capture[7:0] <= 8'd13) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_4 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd0) &&(input_capture[7:0] <= 8'd15) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_5 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd0) &&(input_capture[7:0] <= 8'd1) && 1'b1) ||
     ((input_capture[7:0] >= 8'd8) &&(input_capture[7:0] <= 8'd9) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_6 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd2) &&(input_capture[7:0] <= 8'd3) && 1'b1) ||
     ((input_capture[7:0] >= 8'd10) &&(input_capture[7:0] <= 8'd11) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_7 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd4) &&(input_capture[7:0] <= 8'd7) && 1'b1) ||
     ((input_capture[7:0] >= 8'd12) &&(input_capture[7:0] <= 8'd15) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_8 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd0) &&(input_capture[7:0] <= 8'd1) && 1'b1) ||
     ((input_capture[7:0] >= 8'd8) &&(input_capture[7:0] <= 8'd9) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_ltl0c0_9 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd2) &&(input_capture[7:0] <= 8'd7) && 1'b1) ||
     ((input_capture[7:0] >= 8'd10) &&(input_capture[7:0] <= 8'd15) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule



module Automata_ltl0c0(input clk,
           input run,
           input reset,
           input [7 : 0] symbols
           
           , output ltl0c0_w_out_2
           , output ltl0c0_w_out_4
           , output ltl0c0_w_out_7
           , output ltl0c0_w_out_9);

wire all_input;
wire start_of_data;

assign all_input = 1'b1;
logic start_of_data;
logic start_of_data_reg;
logic start_of_data_reg_ne;

always_ff @ (posedge clk) begin
    if (reset) begin
        start_of_data_reg <= 1;
    end
    else begin
        start_of_data_reg <= 0;
    end
end

always_ff @ (negedge clk) begin
    if (reset) begin
        start_of_data_reg_ne <= 1;
    end
    else begin
        start_of_data_reg_ne <= 0;
    end
end
assign start_of_data = start_of_data_reg & start_of_data_reg_ne & ~reset;




/*wire ltl0c0_w_out_1;
*/

wire ltl0c0_lut_match_1;
wire ltl0c0_w_match_1;

    
    
    

LUT_Match_ltl0c0_1 #(8) lut_match_ltl0c0_1(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_1));


assign ltl0c0_w_match_1 = ltl0c0_lut_match_1 ;

STE #(.fan_in(2),.START_TYPE(1)) ltl0c0_ste_1 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ start_of_data, ltl0c0_w_out_1 }),
                .match(ltl0c0_w_match_1) ,
                .active_state(ltl0c0_w_out_1));




/**/

wire ltl0c0_lut_match_2;
wire ltl0c0_w_match_2;

    
    
    

LUT_Match_ltl0c0_2 #(8) lut_match_ltl0c0_2(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_2));


assign ltl0c0_w_match_2 = ltl0c0_lut_match_2 ;

STE #(.fan_in(2),.START_TYPE(1)) ltl0c0_ste_2 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ start_of_data, ltl0c0_w_out_1 }),
                .match(ltl0c0_w_match_2) ,
                .active_state(ltl0c0_w_out_2));




/*wire ltl0c0_w_out_3;
*/

wire ltl0c0_lut_match_3;
wire ltl0c0_w_match_3;

    
    
    

LUT_Match_ltl0c0_3 #(8) lut_match_ltl0c0_3(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_3));


assign ltl0c0_w_match_3 = ltl0c0_lut_match_3 ;

STE #(.fan_in(2),.START_TYPE(1)) ltl0c0_ste_3 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ start_of_data, ltl0c0_w_out_1 }),
                .match(ltl0c0_w_match_3) ,
                .active_state(ltl0c0_w_out_3));




/**/

wire ltl0c0_lut_match_4;
wire ltl0c0_w_match_4;

    
    
    

LUT_Match_ltl0c0_4 #(8) lut_match_ltl0c0_4(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_4));


assign ltl0c0_w_match_4 = ltl0c0_lut_match_4 ;

STE #(.fan_in(4)) ltl0c0_ste_4 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ ltl0c0_w_out_9, ltl0c0_w_out_2, ltl0c0_w_out_4, ltl0c0_w_out_7 }),
                .match(ltl0c0_w_match_4) ,
                .active_state(ltl0c0_w_out_4));




/*wire ltl0c0_w_out_5;
*/

wire ltl0c0_lut_match_5;
wire ltl0c0_w_match_5;

    
    
    

LUT_Match_ltl0c0_5 #(8) lut_match_ltl0c0_5(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_5));


assign ltl0c0_w_match_5 = ltl0c0_lut_match_5 ;

STE #(.fan_in(2)) ltl0c0_ste_5 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ ltl0c0_w_out_3, ltl0c0_w_out_5 }),
                .match(ltl0c0_w_match_5) ,
                .active_state(ltl0c0_w_out_5));




/*wire ltl0c0_w_out_6;
*/

wire ltl0c0_lut_match_6;
wire ltl0c0_w_match_6;

    
    
    

LUT_Match_ltl0c0_6 #(8) lut_match_ltl0c0_6(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_6));


assign ltl0c0_w_match_6 = ltl0c0_lut_match_6 ;

STE #(.fan_in(2)) ltl0c0_ste_6 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ ltl0c0_w_out_3, ltl0c0_w_out_5 }),
                .match(ltl0c0_w_match_6) ,
                .active_state(ltl0c0_w_out_6));




/**/

wire ltl0c0_lut_match_7;
wire ltl0c0_w_match_7;

    
    
    

LUT_Match_ltl0c0_7 #(8) lut_match_ltl0c0_7(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_7));


assign ltl0c0_w_match_7 = ltl0c0_lut_match_7 ;

STE #(.fan_in(2)) ltl0c0_ste_7 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ ltl0c0_w_out_3, ltl0c0_w_out_5 }),
                .match(ltl0c0_w_match_7) ,
                .active_state(ltl0c0_w_out_7));




/*wire ltl0c0_w_out_8;
*/

wire ltl0c0_lut_match_8;
wire ltl0c0_w_match_8;

    
    
    

LUT_Match_ltl0c0_8 #(8) lut_match_ltl0c0_8(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_8));


assign ltl0c0_w_match_8 = ltl0c0_lut_match_8 ;

STE #(.fan_in(2)) ltl0c0_ste_8 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ ltl0c0_w_out_8, ltl0c0_w_out_6 }),
                .match(ltl0c0_w_match_8) ,
                .active_state(ltl0c0_w_out_8));




/**/

wire ltl0c0_lut_match_9;
wire ltl0c0_w_match_9;

    
    
    

LUT_Match_ltl0c0_9 #(8) lut_match_ltl0c0_9(
                .clk(clk),
                .symbols(symbols),
                .match(ltl0c0_lut_match_9));


assign ltl0c0_w_match_9 = ltl0c0_lut_match_9 ;

STE #(.fan_in(2)) ltl0c0_ste_9 (
                .clk(clk),
                .run(run),
                .reset(reset),
		.start_of_data,
                .income_edges({ ltl0c0_w_out_8, ltl0c0_w_out_6 }),
                .match(ltl0c0_w_match_9) ,
                .active_state(ltl0c0_w_out_9));




endmodule

