

module Top_ModuleC6lw(
                  input clk,
                  input reset,
                  input run,
                  input [7 : 0] symbols
                   , output wire ltl1c6lw
                   , output wire ltl8c6lw
                   , output wire ltl2c6lw
                   , output wire ltl3c6lw
                   , output wire ltl9c6lw
                   , output wire ltl6c6lw
                   , output wire ltl4c6lw
                   , output wire ltl5c6lw
                   , output wire ltl7c6lw
                   , output wire ltl0c6lw
                  
                  );
  wire ltl1c6lw_w_out_4;
  wire ltl1c6lw_w_out_6;
  wire ltl1c6lw_w_out_9;
  wire ltl1c6lw_w_out_11;
  wire ltl8c6lw_w_out_4;
  wire ltl8c6lw_w_out_6;
  wire ltl8c6lw_w_out_9;
  wire ltl8c6lw_w_out_11;
  wire ltl2c6lw_w_out_4;
  wire ltl2c6lw_w_out_6;
  wire ltl2c6lw_w_out_9;
  wire ltl2c6lw_w_out_11;
  wire ltl3c6lw_w_out_4;
  wire ltl3c6lw_w_out_6;
  wire ltl3c6lw_w_out_9;
  wire ltl3c6lw_w_out_11;
  wire ltl9c6lw_w_out_4;
  wire ltl9c6lw_w_out_6;
  wire ltl9c6lw_w_out_9;
  wire ltl9c6lw_w_out_11;
  wire ltl6c6lw_w_out_4;
  wire ltl6c6lw_w_out_6;
  wire ltl6c6lw_w_out_9;
  wire ltl6c6lw_w_out_11;
  wire ltl4c6lw_w_out_4;
  wire ltl4c6lw_w_out_6;
  wire ltl4c6lw_w_out_9;
  wire ltl4c6lw_w_out_11;
  wire ltl5c6lw_w_out_4;
  wire ltl5c6lw_w_out_6;
  wire ltl5c6lw_w_out_9;
  wire ltl5c6lw_w_out_11;
  wire ltl7c6lw_w_out_4;
  wire ltl7c6lw_w_out_6;
  wire ltl7c6lw_w_out_9;
  wire ltl7c6lw_w_out_11;
  wire ltl0c6lw_w_out_4;
  wire ltl0c6lw_w_out_6;
  wire ltl0c6lw_w_out_9;
  wire ltl0c6lw_w_out_11;

assign ltl1c6lw =
  ltl1c6lw_w_out_4 |
  ltl1c6lw_w_out_6 |
  ltl1c6lw_w_out_9 |
  ltl1c6lw_w_out_11 |
1'b0;
assign ltl8c6lw =
  ltl8c6lw_w_out_4 |
  ltl8c6lw_w_out_6 |
  ltl8c6lw_w_out_9 |
  ltl8c6lw_w_out_11 |
1'b0;
assign ltl2c6lw =
  ltl2c6lw_w_out_4 |
  ltl2c6lw_w_out_6 |
  ltl2c6lw_w_out_9 |
  ltl2c6lw_w_out_11 |
1'b0;
assign ltl3c6lw =
  ltl3c6lw_w_out_4 |
  ltl3c6lw_w_out_6 |
  ltl3c6lw_w_out_9 |
  ltl3c6lw_w_out_11 |
1'b0;
assign ltl9c6lw =
  ltl9c6lw_w_out_4 |
  ltl9c6lw_w_out_6 |
  ltl9c6lw_w_out_9 |
  ltl9c6lw_w_out_11 |
1'b0;
assign ltl6c6lw =
  ltl6c6lw_w_out_4 |
  ltl6c6lw_w_out_6 |
  ltl6c6lw_w_out_9 |
  ltl6c6lw_w_out_11 |
1'b0;
assign ltl4c6lw =
  ltl4c6lw_w_out_4 |
  ltl4c6lw_w_out_6 |
  ltl4c6lw_w_out_9 |
  ltl4c6lw_w_out_11 |
1'b0;
assign ltl5c6lw =
  ltl5c6lw_w_out_4 |
  ltl5c6lw_w_out_6 |
  ltl5c6lw_w_out_9 |
  ltl5c6lw_w_out_11 |
1'b0;
assign ltl7c6lw =
  ltl7c6lw_w_out_4 |
  ltl7c6lw_w_out_6 |
  ltl7c6lw_w_out_9 |
  ltl7c6lw_w_out_11 |
1'b0;
assign ltl0c6lw =
  ltl0c6lw_w_out_4 |
  ltl0c6lw_w_out_6 |
  ltl0c6lw_w_out_9 |
  ltl0c6lw_w_out_11 |
1'b0;





Automata_Stage0C6lw automata_stage0(.clk(clk),
                                             .run(run),
                                             .reset(reset),
                                             .top_symbols( symbols ),
                                              .ltl1c6lw_w_out_4(ltl1c6lw_w_out_4),
                                              .ltl1c6lw_w_out_6(ltl1c6lw_w_out_6),
                                              .ltl1c6lw_w_out_9(ltl1c6lw_w_out_9),
                                              .ltl1c6lw_w_out_11(ltl1c6lw_w_out_11),
                                             
                                              .ltl8c6lw_w_out_4(ltl8c6lw_w_out_4),
                                              .ltl8c6lw_w_out_6(ltl8c6lw_w_out_6),
                                              .ltl8c6lw_w_out_9(ltl8c6lw_w_out_9),
                                              .ltl8c6lw_w_out_11(ltl8c6lw_w_out_11),
                                             
                                              .ltl2c6lw_w_out_4(ltl2c6lw_w_out_4),
                                              .ltl2c6lw_w_out_6(ltl2c6lw_w_out_6),
                                              .ltl2c6lw_w_out_9(ltl2c6lw_w_out_9),
                                              .ltl2c6lw_w_out_11(ltl2c6lw_w_out_11),
                                             
                                              .ltl3c6lw_w_out_4(ltl3c6lw_w_out_4),
                                              .ltl3c6lw_w_out_6(ltl3c6lw_w_out_6),
                                              .ltl3c6lw_w_out_9(ltl3c6lw_w_out_9),
                                              .ltl3c6lw_w_out_11(ltl3c6lw_w_out_11),
                                             
                                              .ltl9c6lw_w_out_4(ltl9c6lw_w_out_4),
                                              .ltl9c6lw_w_out_6(ltl9c6lw_w_out_6),
                                              .ltl9c6lw_w_out_9(ltl9c6lw_w_out_9),
                                              .ltl9c6lw_w_out_11(ltl9c6lw_w_out_11),
                                             
                                              .ltl6c6lw_w_out_4(ltl6c6lw_w_out_4),
                                              .ltl6c6lw_w_out_6(ltl6c6lw_w_out_6),
                                              .ltl6c6lw_w_out_9(ltl6c6lw_w_out_9),
                                              .ltl6c6lw_w_out_11(ltl6c6lw_w_out_11),
                                             
                                              .ltl4c6lw_w_out_4(ltl4c6lw_w_out_4),
                                              .ltl4c6lw_w_out_6(ltl4c6lw_w_out_6),
                                              .ltl4c6lw_w_out_9(ltl4c6lw_w_out_9),
                                              .ltl4c6lw_w_out_11(ltl4c6lw_w_out_11),
                                             
                                              .ltl5c6lw_w_out_4(ltl5c6lw_w_out_4),
                                              .ltl5c6lw_w_out_6(ltl5c6lw_w_out_6),
                                              .ltl5c6lw_w_out_9(ltl5c6lw_w_out_9),
                                              .ltl5c6lw_w_out_11(ltl5c6lw_w_out_11),
                                             
                                              .ltl7c6lw_w_out_4(ltl7c6lw_w_out_4),
                                              .ltl7c6lw_w_out_6(ltl7c6lw_w_out_6),
                                              .ltl7c6lw_w_out_9(ltl7c6lw_w_out_9),
                                              .ltl7c6lw_w_out_11(ltl7c6lw_w_out_11),
                                             
                                              .ltl0c6lw_w_out_4(ltl0c6lw_w_out_4),
                                              .ltl0c6lw_w_out_6(ltl0c6lw_w_out_6),
                                              .ltl0c6lw_w_out_9(ltl0c6lw_w_out_9),
                                              .ltl0c6lw_w_out_11(ltl0c6lw_w_out_11),
                                             
                                             .out_symbols(),
                                             .out_reset()
                                             );




endmodule
