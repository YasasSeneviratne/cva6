





/*
******************** Summary {}********************
total nodes = 121
total reports = 44
total edges = 242
average symbols len = 12.8347107438
#######################################################
*/

module Automata_Stage0C0(input clk,
                    input run,
                    input reset,
                    input [7 : 0] top_symbols
                    , output ltl2c0_w_out_4
                    , output ltl2c0_w_out_6
                    , output ltl2c0_w_out_9
                    , output ltl2c0_w_out_11
                    
                    , output ltl9c0_w_out_4
                    , output ltl9c0_w_out_6
                    , output ltl9c0_w_out_9
                    , output ltl9c0_w_out_11
                    
                    , output ltl0c0_w_out_4
                    , output ltl0c0_w_out_6
                    , output ltl0c0_w_out_9
                    , output ltl0c0_w_out_11
                    
                    , output ltl8c0_w_out_4
                    , output ltl8c0_w_out_6
                    , output ltl8c0_w_out_9
                    , output ltl8c0_w_out_11
                    
                    , output ltl1c0_w_out_4
                    , output ltl1c0_w_out_6
                    , output ltl1c0_w_out_9
                    , output ltl1c0_w_out_11
                    
                    , output ltl4c0_w_out_4
                    , output ltl4c0_w_out_6
                    , output ltl4c0_w_out_9
                    , output ltl4c0_w_out_11
                    
                    , output ltl3c0_w_out_4
                    , output ltl3c0_w_out_6
                    , output ltl3c0_w_out_9
                    , output ltl3c0_w_out_11
                    
                    , output ltl10c0_w_out_4
                    , output ltl10c0_w_out_6
                    , output ltl10c0_w_out_9
                    , output ltl10c0_w_out_11
                    
                    , output ltl7c0_w_out_4
                    , output ltl7c0_w_out_6
                    , output ltl7c0_w_out_9
                    , output ltl7c0_w_out_11
                    
                    , output ltl5c0_w_out_4
                    , output ltl5c0_w_out_6
                    , output ltl5c0_w_out_9
                    , output ltl5c0_w_out_11
                    
                    , output ltl6c0_w_out_4
                    , output ltl6c0_w_out_6
                    , output ltl6c0_w_out_9
                    , output ltl6c0_w_out_11
                    ,
                    output reg[7 : 0] out_symbols,
                    output reg out_reset
                    );

always @(posedge clk)
begin
    if (run == 1)
        out_symbols <= top_symbols;
        out_reset <= reset;
end



Automata_ltl2c0 automata_ltl2c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl2c0_w_out_4(ltl2c0_w_out_4)
                        , .ltl2c0_w_out_6(ltl2c0_w_out_6)
                        , .ltl2c0_w_out_9(ltl2c0_w_out_9)
                        , .ltl2c0_w_out_11(ltl2c0_w_out_11)
                    );

Automata_ltl9c0 automata_ltl9c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl9c0_w_out_4(ltl9c0_w_out_4)
                        , .ltl9c0_w_out_6(ltl9c0_w_out_6)
                        , .ltl9c0_w_out_9(ltl9c0_w_out_9)
                        , .ltl9c0_w_out_11(ltl9c0_w_out_11)
                    );

Automata_ltl0c0 automata_ltl0c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl0c0_w_out_4(ltl0c0_w_out_4)
                        , .ltl0c0_w_out_6(ltl0c0_w_out_6)
                        , .ltl0c0_w_out_9(ltl0c0_w_out_9)
                        , .ltl0c0_w_out_11(ltl0c0_w_out_11)
                    );

Automata_ltl8c0 automata_ltl8c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl8c0_w_out_4(ltl8c0_w_out_4)
                        , .ltl8c0_w_out_6(ltl8c0_w_out_6)
                        , .ltl8c0_w_out_9(ltl8c0_w_out_9)
                        , .ltl8c0_w_out_11(ltl8c0_w_out_11)
                    );

Automata_ltl1c0 automata_ltl1c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl1c0_w_out_4(ltl1c0_w_out_4)
                        , .ltl1c0_w_out_6(ltl1c0_w_out_6)
                        , .ltl1c0_w_out_9(ltl1c0_w_out_9)
                        , .ltl1c0_w_out_11(ltl1c0_w_out_11)
                    );

Automata_ltl4c0 automata_ltl4c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl4c0_w_out_4(ltl4c0_w_out_4)
                        , .ltl4c0_w_out_6(ltl4c0_w_out_6)
                        , .ltl4c0_w_out_9(ltl4c0_w_out_9)
                        , .ltl4c0_w_out_11(ltl4c0_w_out_11)
                    );

Automata_ltl3c0 automata_ltl3c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl3c0_w_out_4(ltl3c0_w_out_4)
                        , .ltl3c0_w_out_6(ltl3c0_w_out_6)
                        , .ltl3c0_w_out_9(ltl3c0_w_out_9)
                        , .ltl3c0_w_out_11(ltl3c0_w_out_11)
                    );

Automata_ltl10c0 automata_ltl10c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl10c0_w_out_4(ltl10c0_w_out_4)
                        , .ltl10c0_w_out_6(ltl10c0_w_out_6)
                        , .ltl10c0_w_out_9(ltl10c0_w_out_9)
                        , .ltl10c0_w_out_11(ltl10c0_w_out_11)
                    );

Automata_ltl7c0 automata_ltl7c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl7c0_w_out_4(ltl7c0_w_out_4)
                        , .ltl7c0_w_out_6(ltl7c0_w_out_6)
                        , .ltl7c0_w_out_9(ltl7c0_w_out_9)
                        , .ltl7c0_w_out_11(ltl7c0_w_out_11)
                    );

Automata_ltl5c0 automata_ltl5c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl5c0_w_out_4(ltl5c0_w_out_4)
                        , .ltl5c0_w_out_6(ltl5c0_w_out_6)
                        , .ltl5c0_w_out_9(ltl5c0_w_out_9)
                        , .ltl5c0_w_out_11(ltl5c0_w_out_11)
                    );

Automata_ltl6c0 automata_ltl6c0 (
                     .clk(clk),
                     .run(run),
                     .reset(reset),
                        .symbols(top_symbols )
                        , .ltl6c0_w_out_4(ltl6c0_w_out_4)
                        , .ltl6c0_w_out_6(ltl6c0_w_out_6)
                        , .ltl6c0_w_out_9(ltl6c0_w_out_9)
                        , .ltl6c0_w_out_11(ltl6c0_w_out_11)
                    );


























    



 










endmodule
