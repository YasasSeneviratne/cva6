

module Top_ModuleC3lw(
                  input clk,
                  input reset,
                  input run,
                  input [7 : 0] symbols
                   , output wire ltl8c3lw
                   , output wire ltl0c3lw
                   , output wire ltl9c3lw
                   , output wire ltl3c3lw
                   , output wire ltl6c3lw
                   , output wire ltl4c3lw
                   , output wire ltl7c3lw
                   , output wire ltl5c3lw
                   , output wire ltl2c3lw
                   , output wire ltl1c3lw
                  
                  );
  wire ltl8c3lw_w_out_4;
  wire ltl8c3lw_w_out_6;
  wire ltl8c3lw_w_out_9;
  wire ltl8c3lw_w_out_11;
  wire ltl0c3lw_w_out_4;
  wire ltl0c3lw_w_out_6;
  wire ltl0c3lw_w_out_9;
  wire ltl0c3lw_w_out_11;
  wire ltl9c3lw_w_out_4;
  wire ltl9c3lw_w_out_6;
  wire ltl9c3lw_w_out_9;
  wire ltl9c3lw_w_out_11;
  wire ltl3c3lw_w_out_4;
  wire ltl3c3lw_w_out_6;
  wire ltl3c3lw_w_out_9;
  wire ltl3c3lw_w_out_11;
  wire ltl6c3lw_w_out_4;
  wire ltl6c3lw_w_out_6;
  wire ltl6c3lw_w_out_9;
  wire ltl6c3lw_w_out_11;
  wire ltl4c3lw_w_out_4;
  wire ltl4c3lw_w_out_6;
  wire ltl4c3lw_w_out_9;
  wire ltl4c3lw_w_out_11;
  wire ltl7c3lw_w_out_4;
  wire ltl7c3lw_w_out_6;
  wire ltl7c3lw_w_out_9;
  wire ltl7c3lw_w_out_11;
  wire ltl5c3lw_w_out_4;
  wire ltl5c3lw_w_out_6;
  wire ltl5c3lw_w_out_9;
  wire ltl5c3lw_w_out_11;
  wire ltl2c3lw_w_out_4;
  wire ltl2c3lw_w_out_6;
  wire ltl2c3lw_w_out_9;
  wire ltl2c3lw_w_out_11;
  wire ltl1c3lw_w_out_4;
  wire ltl1c3lw_w_out_6;
  wire ltl1c3lw_w_out_9;
  wire ltl1c3lw_w_out_11;

assign ltl8c3lw =
  ltl8c3lw_w_out_4 |
  ltl8c3lw_w_out_6 |
  ltl8c3lw_w_out_9 |
  ltl8c3lw_w_out_11 |
1'b0;
assign ltl0c3lw =
  ltl0c3lw_w_out_4 |
  ltl0c3lw_w_out_6 |
  ltl0c3lw_w_out_9 |
  ltl0c3lw_w_out_11 |
1'b0;
assign ltl9c3lw =
  ltl9c3lw_w_out_4 |
  ltl9c3lw_w_out_6 |
  ltl9c3lw_w_out_9 |
  ltl9c3lw_w_out_11 |
1'b0;
assign ltl3c3lw =
  ltl3c3lw_w_out_4 |
  ltl3c3lw_w_out_6 |
  ltl3c3lw_w_out_9 |
  ltl3c3lw_w_out_11 |
1'b0;
assign ltl6c3lw =
  ltl6c3lw_w_out_4 |
  ltl6c3lw_w_out_6 |
  ltl6c3lw_w_out_9 |
  ltl6c3lw_w_out_11 |
1'b0;
assign ltl4c3lw =
  ltl4c3lw_w_out_4 |
  ltl4c3lw_w_out_6 |
  ltl4c3lw_w_out_9 |
  ltl4c3lw_w_out_11 |
1'b0;
assign ltl7c3lw =
  ltl7c3lw_w_out_4 |
  ltl7c3lw_w_out_6 |
  ltl7c3lw_w_out_9 |
  ltl7c3lw_w_out_11 |
1'b0;
assign ltl5c3lw =
  ltl5c3lw_w_out_4 |
  ltl5c3lw_w_out_6 |
  ltl5c3lw_w_out_9 |
  ltl5c3lw_w_out_11 |
1'b0;
assign ltl2c3lw =
  ltl2c3lw_w_out_4 |
  ltl2c3lw_w_out_6 |
  ltl2c3lw_w_out_9 |
  ltl2c3lw_w_out_11 |
1'b0;
assign ltl1c3lw =
  ltl1c3lw_w_out_4 |
  ltl1c3lw_w_out_6 |
  ltl1c3lw_w_out_9 |
  ltl1c3lw_w_out_11 |
1'b0;





Automata_Stage0C3lw automata_stage0(.clk(clk),
                                             .run(run),
                                             .reset(reset),
                                             .top_symbols( symbols ),
                                              .ltl8c3lw_w_out_4(ltl8c3lw_w_out_4),
                                              .ltl8c3lw_w_out_6(ltl8c3lw_w_out_6),
                                              .ltl8c3lw_w_out_9(ltl8c3lw_w_out_9),
                                              .ltl8c3lw_w_out_11(ltl8c3lw_w_out_11),
                                             
                                              .ltl0c3lw_w_out_4(ltl0c3lw_w_out_4),
                                              .ltl0c3lw_w_out_6(ltl0c3lw_w_out_6),
                                              .ltl0c3lw_w_out_9(ltl0c3lw_w_out_9),
                                              .ltl0c3lw_w_out_11(ltl0c3lw_w_out_11),
                                             
                                              .ltl9c3lw_w_out_4(ltl9c3lw_w_out_4),
                                              .ltl9c3lw_w_out_6(ltl9c3lw_w_out_6),
                                              .ltl9c3lw_w_out_9(ltl9c3lw_w_out_9),
                                              .ltl9c3lw_w_out_11(ltl9c3lw_w_out_11),
                                             
                                              .ltl3c3lw_w_out_4(ltl3c3lw_w_out_4),
                                              .ltl3c3lw_w_out_6(ltl3c3lw_w_out_6),
                                              .ltl3c3lw_w_out_9(ltl3c3lw_w_out_9),
                                              .ltl3c3lw_w_out_11(ltl3c3lw_w_out_11),
                                             
                                              .ltl6c3lw_w_out_4(ltl6c3lw_w_out_4),
                                              .ltl6c3lw_w_out_6(ltl6c3lw_w_out_6),
                                              .ltl6c3lw_w_out_9(ltl6c3lw_w_out_9),
                                              .ltl6c3lw_w_out_11(ltl6c3lw_w_out_11),
                                             
                                              .ltl4c3lw_w_out_4(ltl4c3lw_w_out_4),
                                              .ltl4c3lw_w_out_6(ltl4c3lw_w_out_6),
                                              .ltl4c3lw_w_out_9(ltl4c3lw_w_out_9),
                                              .ltl4c3lw_w_out_11(ltl4c3lw_w_out_11),
                                             
                                              .ltl7c3lw_w_out_4(ltl7c3lw_w_out_4),
                                              .ltl7c3lw_w_out_6(ltl7c3lw_w_out_6),
                                              .ltl7c3lw_w_out_9(ltl7c3lw_w_out_9),
                                              .ltl7c3lw_w_out_11(ltl7c3lw_w_out_11),
                                             
                                              .ltl5c3lw_w_out_4(ltl5c3lw_w_out_4),
                                              .ltl5c3lw_w_out_6(ltl5c3lw_w_out_6),
                                              .ltl5c3lw_w_out_9(ltl5c3lw_w_out_9),
                                              .ltl5c3lw_w_out_11(ltl5c3lw_w_out_11),
                                             
                                              .ltl2c3lw_w_out_4(ltl2c3lw_w_out_4),
                                              .ltl2c3lw_w_out_6(ltl2c3lw_w_out_6),
                                              .ltl2c3lw_w_out_9(ltl2c3lw_w_out_9),
                                              .ltl2c3lw_w_out_11(ltl2c3lw_w_out_11),
                                             
                                              .ltl1c3lw_w_out_4(ltl1c3lw_w_out_4),
                                              .ltl1c3lw_w_out_6(ltl1c3lw_w_out_6),
                                              .ltl1c3lw_w_out_9(ltl1c3lw_w_out_9),
                                              .ltl1c3lw_w_out_11(ltl1c3lw_w_out_11),
                                             
                                             .out_symbols(),
                                             .out_reset()
                                             );




endmodule
